Begin3
Language:    SV, 850, Swedish
Title:       cabextract
Description: cabextract kan extrahera filer fr�n en m�ngd olika Microsoft CAB-format.
Keywords:    cab, komprimerat, arkiv
End
